module Mux(input [5:0]num,output reg [13:0]disp);
always@(*)
case(num)
6'd00: disp = 14'b1111110_1111110;
6'd01: disp = 14'b1111110_0110000;
6'd02: disp = 14'b1111110_1101101;
6'd03: disp = 14'b1111110_1111001;
6'd04: disp = 14'b1111110_0010011;
6'd05: disp = 14'b1111110_0011011;
6'd06: disp = 14'b1111110_1011111;
6'd07: disp = 14'b1111110_1110000;
6'd08: disp = 14'b1111110_1111111;
6'd09: disp = 14'b1111110_1111011;
6'd10: disp = 14'b0110000_1111110;
6'd11: disp = 14'b0110000_0110000;
6'd12: disp = 14'b0110000_1101101;
6'd13: disp = 14'b0110000_1111001;
6'd14: disp = 14'b0110000_0010011;
6'd15: disp = 14'b0110000_0011011;
6'd16: disp = 14'b0110000_1011111;
6'd17: disp = 14'b0110000_1110000;
6'd18: disp = 14'b0110000_1111111;
6'd19: disp = 14'b0110000_1111011;
6'd20: disp = 14'b1101101_1111110;
6'd21: disp = 14'b1101101_0110000;
6'd22: disp = 14'b1101101_1101101;
6'd23: disp = 14'b1101101_1111001;
6'd24: disp = 14'b1101101_0010011;
6'd25: disp = 14'b1101101_0011011;
6'd26: disp = 14'b1101101_1011111;
6'd27: disp = 14'b1101101_1110000;
6'd28: disp = 14'b1101101_1111111;
6'd29: disp = 14'b1101101_1111011;
6'd30: disp = 14'b1111001_1111110;
6'd31: disp = 14'b1111001_0110000;
6'd32: disp = 14'b1111001_1101101;
6'd33: disp = 14'b1111001_1111001;
6'd34: disp = 14'b1111001_0010011;
6'd35: disp = 14'b1111001_0011011;
6'd36: disp = 14'b1111001_1011111;
6'd37: disp = 14'b1111001_1110000;
6'd38: disp = 14'b1111001_1111111;
6'd39: disp = 14'b1111001_1111011;
6'd40: disp = 14'b0010011_1111110;
6'd41: disp = 14'b0010011_0110000;
6'd42: disp = 14'b0010011_1101101;
6'd43: disp = 14'b0010011_1111001;
6'd44: disp = 14'b0010011_0010011;
6'd45: disp = 14'b0010011_0011011;
6'd46: disp = 14'b0010011_1011111;
6'd47: disp = 14'b0010011_1110000;
6'd48: disp = 14'b0010011_1111111;
6'd49: disp = 14'b0010011_1111011;
6'd50: disp = 14'b0011011_1111110;
6'd51: disp = 14'b0011011_0110000;
6'd52: disp = 14'b0011011_1101101;
6'd53: disp = 14'b0011011_1111001;
6'd54: disp = 14'b0011011_0010011;
6'd55: disp = 14'b0011011_0011011;
6'd56: disp = 14'b0011011_1011111;
6'd57: disp = 14'b0011011_1110000;
6'd58: disp = 14'b0011011_1111111;
6'd59: disp = 14'b0011011_1111011;
endcase
endmodule
